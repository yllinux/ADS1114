library verilog;
use verilog.vl_types.all;
entity SEG7_TOP_vlg_tst is
end SEG7_TOP_vlg_tst;
